module segled(
    input  wire [3:0] x,
    output wire [6:0] z
);

assign z = (x == 0) ? 7'b1000000 :
			(x == 1) ? 7'b1111001 :
			(x == 2) ? 7'b0100100 :
			(x == 3) ? 7'b0110000 :
			(x == 4) ? 7'b0011001 :
			(x == 5) ? 7'b0010010 :
			(x == 6) ? 7'b0000010 :
			(x == 7) ? 7'b1111000 :
			(x == 8) ? 7'b0000000 :
			(x == 9) ? 7'b0010000 :
			(x == 10)? 7'b0001000 :
			(x == 11)? 7'b0000011 :
			(x == 12)? 7'b1000110 :
			(x == 13)? 7'b0100001 :
			(x == 14)? 7'b0000110 :
			7'b0001110;
endmodule
